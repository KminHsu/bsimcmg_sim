
* .options output initial_interval=5e-6
* .options timeint reltol=1e-6 abstol=1e-6 method=trap maxord=1
* * V1 1 0 dc 1.0
* *V1 1 0 1 AC 1 PULSE 1 0 500m 1000m
* *V1 1 0 1 AC 1 PULSE 1 0 1000m 0m 2000m
* V1 1 0 PULSE 1 0 50m 0m 100m
* R1 1 2 1
* C1 2 0 1
* *.op
* *.ic V(2)=0.5
* .tran 0n 100m
* .print tran format=csv v(*) 

*.OPTIONS LIST NODE POST
.options output initial_interval=1e-8
.options timeint reltol=1e-6 abstol=1e-6 method=trap maxord=1
*.OP
.TRAN 0 2U
.PRINT TRAN format=csv PRECISION=20 V(1) V(2) I(R2) I(C1)
*V1 1 0 10 AC 1 PULSE 0 5 10N 20N 20N 500N 2U
V1 1 0 10 AC 1 PULSE 0 5 0 0 0 5e-7 2U
R1 1 2 1K
R2 2 0 1K
C1 2 0 .001U
.END


